`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:2**8-1];

    initial begin
        $readmemh("code.mem", rom);


        //rom[x]=32'b fucn7 _ rs2 _ rs1 _f3 _ rd  _ op // R-Type
        //rom[0] = 32'b0000000_00001_00010_000_00100_0110011;  // add x4, x2, x1 : regfile 4번주소 = 12+11 = 23
        //rom[1] = 32'b0100000_00001_00010_000_00101_0110011;  // sub x5, x2, x1 : 5번 주소 = 12-11 = 1
        //rom[2] = 32'b0000000_00000_00011_111_00110_0110011;  // and x6, x3, x0 : 6번 주소 = 13 and 0 = 0
        //rom[3] = 32'b0000000_00000_00011_110_00111_0110011;  // or  x7, x3, x0 : 7번 주소 = 13 or 0 = 13
        //rom[4] = 32'b0000000_00010_00011_100_01000_0110011;  // xor x8, x3, x2 : 8번 주소 = 00001 = 1

        //rom[5] = 32'b0000000_11110_00001_001_01001_0110011;  // sll x9, x1, x30 : 9번 주소 = 11<<1 = 01011<<1 = 10110: 22 
        //rom[6] = 32'b0000000_11110_01110_101_01010_0110011;  // srl x10, x14, x30 : 10번 주소 = 위의 x9 값 >> 1 = 1011 (11)
        //rom[7] = 32'b0100000_11110_11111_101_01011_0110011; // sra x11, x31, x30 : 11번 주소 = -2 >>> 1 : _1110(_FFFE) >>> 1 = _1111(_FFFF)
        //rom[8] = 32'b0000000_00000_11111_010_01100_0110011; // slt x12, x31, x0 : 12번 주소는 x0(0) < x1(11) 이면 1
        //rom[9] = 32'b0000000_00000_00001_011_01101_0110011; // sltu x13, x1, x0 : 13번 주소 = x1(11) < x0(0) 이므로 0이고 0-extend

        //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // S-Type
        //rom[5] = 32'b0000000_00001_00000_000_01100_0100011; // sb x1, 12(x0) : RAM(addr[12] = mem[3])에 rs2(11) 8bit 쓰기 
        //rom[6] = 32'b0000000_00011_00000_001_10000_0100011; // sh x3, 4(x0)  :RAM(addr[16] = mem[4])에 rs2(13) 16bit 쓰기
        //rom[7] = 32'b0000000_00010_00000_010_01000_0100011;  // sw x2, 8(x0) : RAM(addr[8] = mem[2])에 rs2(12) 32bit 쓰기
        

        //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // B-Type
        //rom[10] = 32'b00000000000100001000010001100011;  // beq x1, x1, 8 : x1 == x1 참이므로 PC += 8 = rom[12] = PC[48]
        //rom[12] = 32'b00000000001000001001010001100011; // bne x1, x2, 8 : x1 != x2 참이므로 PC += 8 = rom[14] = PC[56] 
        //rom[14] = 32'b00000000001011111100010001100011; // blt x31, x2, 8 : x31 < x2 참이므로 PC += 8 = rom[16] = PC[64]
        //rom[16] = 32'b00000001111100010101010001100011; // bge x2, x31, 8 : x2 >= x31 참 PC += 8 = rom[18] = PC[72]
        //rom[18] = 32'b00000000001000001110010001100011; // bltu x1, x2, 8 : x1 < x2 참이므로 rom[20] = PC[80]
        //rom[20] = 32'b00000010000100010111010001100011; // bgeu x2, x1, 40 : x2 >= x1 참이므로 rom[30] = PC[120] = 1(regfile)

        //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // L-Type
        //rom[5] = 32'b00000000100000000000010100000011; // lb x10, 8(x0) : RAM의 2번 주소에서 값을 꺼내와 RegFile의 10번 주소에 쓰기 : 2를 singed extend 해서 쓰기 : 2
        //rom[6] = 32'b00000000110000000001010110000011; // lh x11, 12(x0) : 3번 주소(4) 를 RegFile의 11번 주소에 쓰기 : 4
        //rom[7] = 32'b00000001000000000010011000000011;  // lw x12, 16(x0) : 4번 주소(8)을 12에 쓸꺼니까 : 8
        //rom[8] = 32'b00000001010000000100011010000011; // lbu x13, 20(x0) : 5번 주소(-2)를 13번에 쓰기 : unsigned로 읽기 : 254
        //rom[9] = 32'b00000001100000000101011100000011; // lhu x14, 24(x0) : 6번 주소(-4)를 14번에 쓰기 : unsigned: 65532

        //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // I-Type
        //rom[10] = 32'b000000000010_00001_000_01110_0010011;  // addi x14, x1, 2 : 11 + 2 = 13
        //rom[11] = 32'b00000000101011111010011110010011;  // slti x15, x31, 10 : -2 < 10 ? -> 1
        //rom[12] = 32'b00000000101000001011100000010011;  // sltiu x16, x1, 10 : 11<10 ? -> 0
        //rom[13] = 32'b00000000101000001100100010010011;  // xori x17, x1, 10 : 11^10 -> 1
        //rom[14] = 32'b00000000101000001110100100010011;  // ori x18, x1, 10 : 11|10 -> 11 (1011)
        //rom[15] = 32'b00000000101000001111100110010011;  // andi x19, x1, 10 : 11 & 10 -> 10 (1010)

        //rom[16] = 32'b00000000001000001001101000010011; // slli x20, x1, 2 : 11 << 2 = 44 (101100)
        //rom[17] = 32'b00000000000100001101101010010011; // srli x21, x1, 1 : 11 >> 1 = 5(101)
        //rom[18] = 32'b01000000000111111101101100010011; // srai x22, x31, 1 : -2 >>> 1 = -1 (...11111)

        //LU-Type
        //rom[10] = 32'b00000000000000000010011100110111;  // lui x14, 2 : RegFile 14번 주소에 2 << 12 = 8192
        //AU-Type
        //rom[11] = 32'b00000000000000000001011110010111; // auipc x15, 1 : 15번 주소 값 = PC(44) + 4048 = 4092

        //J-Type
        //rom[10] = 32'b00000000100000000000011101101111; // jal x14, 8 : regfile 14번에 40+4 = 44, PC = 40 + 8 = 48
        //JL-Type
        //rom[12] = 32'b00000000100000000000011111100111; // jalr x15, 8(x0) : regfile 15번에 48+4 = 52, PC = x0(0) + 8 = 56
    
    end

    assign data = rom[addr[31:2]];
endmodule
